//
// Copyright (c) 2015 University of Cambridge
// All rights reserved.
//
//
//  File:
//        output_port_lookup_cpu_regs.v
//
//  Module:
//        output_port_lookup_cpu_regs
//
//  Description:
//        This file is automatically generated with the registers towards the CPU/Software
//
// This software was developed by Stanford University and the University of Cambridge Computer Laboratory
// under National Science Foundation under Grant No. CNS-0855268,
// the University of Cambridge Computer Laboratory under EPSRC INTERNET Project EP/H040536/1 and
// by the University of Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-11-C-0249 ("MRC2"),
// as part of the DARPA MRC research programme.
//
// @NETFPGA_LICENSE_HEADER_START@
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//  http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
// @NETFPGA_LICENSE_HEADER_END@
//

`include "output_port_lookup_cpu_regs_defines.v"
module output_port_lookup_cpu_regs #
(
parameter C_BASE_ADDRESS        = 32'h00000000,
parameter C_S_AXI_DATA_WIDTH    = 32,
parameter C_S_AXI_ADDR_WIDTH    = 32
)
(
    // General ports
    input       clk,
    input       resetn,
    // Global Registers
    input       cpu_resetn_soft,
    output reg  resetn_soft,
    output reg  resetn_sync,

   // Register ports
    input      [`REG_ID_BITS]    id_reg,
    input      [`REG_VERSION_BITS]    version_reg,
    output reg [`REG_RESET_BITS]    reset_reg,
    input      [`REG_FLIP_BITS]    ip2cpu_flip_reg,
    output reg [`REG_FLIP_BITS]    cpu2ip_flip_reg,
    input      [`REG_DEBUG_BITS]    ip2cpu_debug_reg,
    output reg [`REG_DEBUG_BITS]    cpu2ip_debug_reg,
    input      [`REG_PKT_SENT_FROM_CPU_CNTR_BITS]    pkt_sent_from_cpu_cntr_reg,
    output reg                          pkt_sent_from_cpu_cntr_reg_clear,
    input      [`REG_PKT_SENT_TO_CPU_OPTIONS_VER_CNTR_BITS]    pkt_sent_to_cpu_options_ver_cntr_reg,
    output reg                          pkt_sent_to_cpu_options_ver_cntr_reg_clear,
    input      [`REG_PKT_SENT_TO_CPU_BAD_TTL_CNTR_BITS]    pkt_sent_to_cpu_bad_ttl_cntr_reg,
    output reg                          pkt_sent_to_cpu_bad_ttl_cntr_reg_clear,
    input      [`REG_PKT_SENT_TO_CPU_DEST_IP_HIT_CNTR_BITS]    pkt_sent_to_cpu_dest_ip_hit_cntr_reg,
    output reg                          pkt_sent_to_cpu_dest_ip_hit_cntr_reg_clear,
    input      [`REG_PKT_FORWARDED_CNTR_BITS]    pkt_forwarded_cntr_reg,
    output reg                          pkt_forwarded_cntr_reg_clear,
    input      [`REG_PKT_DROPPED_CHECKSUM_CNTR_BITS]    pkt_dropped_checksum_cntr_reg,
    output reg                          pkt_dropped_checksum_cntr_reg_clear,
    input      [`REG_PKT_SENT_TO_CPU_NON_IP_CNTR_BITS]    pkt_sent_to_cpu_non_ip_cntr_reg,
    output reg                          pkt_sent_to_cpu_non_ip_cntr_reg_clear,
    input      [`REG_PKT_SENT_TO_CPU_ARP_MISS_CNTR_BITS]    pkt_sent_to_cpu_arp_miss_cntr_reg,
    output reg                          pkt_sent_to_cpu_arp_miss_cntr_reg_clear,
    input      [`REG_PKT_SENT_TO_CPU_LPM_MISS_CNTR_BITS]    pkt_sent_to_cpu_lpm_miss_cntr_reg,
    output reg                          pkt_sent_to_cpu_lpm_miss_cntr_reg_clear,
    input      [`REG_PKT_DROPPED_WRONG_DST_MAC_CNTR_BITS]    pkt_dropped_wrong_dst_mac_cntr_reg,
    output reg                          pkt_dropped_wrong_dst_mac_cntr_reg_clear,
    output reg [`REG_MAC_0_HI_BITS]    mac_0_hi_reg,
    output reg [`REG_MAC_0_LOW_BITS]    mac_0_low_reg,
    output reg [`REG_MAC_1_HI_BITS]    mac_1_hi_reg,
    output reg [`REG_MAC_1_LOW_BITS]    mac_1_low_reg,
    output reg [`REG_MAC_2_HI_BITS]    mac_2_hi_reg,
    output reg [`REG_MAC_2_LOW_BITS]    mac_2_low_reg,
    output reg [`REG_MAC_3_HI_BITS]    mac_3_hi_reg,
    output reg [`REG_MAC_3_LOW_BITS]    mac_3_low_reg,
    output  reg [`MEM_IP_LPM_TCAM_ADDR_BITS]    ip_lpm_tcam_addr,
    output  reg [127:0]    ip_lpm_tcam_data,
    output  reg                         ip_lpm_tcam_rd_wrn,
    output  reg                         ip_lpm_tcam_cmd_valid,
    input       [127:0]    ip_lpm_tcam_reply,
    input                               ip_lpm_tcam_reply_valid,
    output  reg [`MEM_IP_ARP_CAM_ADDR_BITS]    ip_arp_cam_addr,
    output  reg [127:0]    ip_arp_cam_data,
    output  reg                         ip_arp_cam_rd_wrn,
    output  reg                         ip_arp_cam_cmd_valid,
    input       [127:0]    ip_arp_cam_reply,
    input                               ip_arp_cam_reply_valid,
    output  reg [`MEM_DEST_IP_CAM_ADDR_BITS]    dest_ip_cam_addr,
    output  reg [127:0]    dest_ip_cam_data,
    output  reg                         dest_ip_cam_rd_wrn,
    output  reg                         dest_ip_cam_cmd_valid,
    input       [127:0]    dest_ip_cam_reply,
    input                               dest_ip_cam_reply_valid,

    // AXI Lite ports
    input                                     S_AXI_ACLK,
    input                                     S_AXI_ARESETN,
    input      [C_S_AXI_ADDR_WIDTH-1 : 0]     S_AXI_AWADDR,
    input                                     S_AXI_AWVALID,
    input      [C_S_AXI_DATA_WIDTH-1 : 0]     S_AXI_WDATA,
    input      [C_S_AXI_DATA_WIDTH/8-1 : 0]   S_AXI_WSTRB,
    input                                     S_AXI_WVALID,
    input                                     S_AXI_BREADY,
    input      [C_S_AXI_ADDR_WIDTH-1 : 0]     S_AXI_ARADDR,
    input                                     S_AXI_ARVALID,
    input                                     S_AXI_RREADY,
    output                                    S_AXI_ARREADY,
    output     [C_S_AXI_DATA_WIDTH-1 : 0]     S_AXI_RDATA,
    output     [1 : 0]                        S_AXI_RRESP,
    output                                    S_AXI_RVALID,
    output                                    S_AXI_WREADY,
    output     [1 :0]                         S_AXI_BRESP,
    output                                    S_AXI_BVALID,
    output                                    S_AXI_AWREADY

);

    // AXI4LITE signals
    reg [C_S_AXI_ADDR_WIDTH-1 : 0]      axi_awaddr;
    reg                                 axi_awready;
    reg                                 axi_wready;
    reg [1 : 0]                         axi_bresp;
    reg                                 axi_bvalid;
    reg [C_S_AXI_ADDR_WIDTH-1 : 0]      axi_araddr;
    reg                                 axi_arready;
    reg [C_S_AXI_DATA_WIDTH-1 : 0]      axi_rdata;
    reg [1 : 0]                         axi_rresp;
    reg                                 axi_rvalid;

    reg                                 resetn_sync_d;
    wire                                reg_rden;
    wire                                reg_wren;
    reg [C_S_AXI_DATA_WIDTH-1:0]        reg_data_out;
    integer                             byte_index;
    reg                                 pkt_sent_from_cpu_cntr_reg_clear_d;
    reg                                 pkt_sent_to_cpu_options_ver_cntr_reg_clear_d;
    reg                                 pkt_sent_to_cpu_bad_ttl_cntr_reg_clear_d;
    reg                                 pkt_sent_to_cpu_dest_ip_hit_cntr_reg_clear_d;
    reg                                 pkt_forwarded_cntr_reg_clear_d;
    reg                                 pkt_dropped_checksum_cntr_reg_clear_d;
    reg                                 pkt_sent_to_cpu_non_ip_cntr_reg_clear_d;
    reg                                 pkt_sent_to_cpu_arp_miss_cntr_reg_clear_d;
    reg                                 pkt_sent_to_cpu_lpm_miss_cntr_reg_clear_d;
    reg                                 pkt_dropped_wrong_dst_mac_cntr_reg_clear_d;
    reg      [`REG_INDIRECTADDRESS_BITS] indirectaddress_reg;
    reg      [`REG_INDIRECTWRDATA_A_HI_BITS] indirectwrdata_a_hi_reg;
    reg      [`REG_INDIRECTWRDATA_A_LOW_BITS] indirectwrdata_a_low_reg;
    reg      [`REG_INDIRECTWRDATA_B_HI_BITS] indirectwrdata_b_hi_reg;
    reg      [`REG_INDIRECTWRDATA_B_LOW_BITS] indirectwrdata_b_low_reg;
    reg      [`REG_INDIRECTREPLY_A_HI_BITS] indirectreply_a_hi_reg;
    reg      [`REG_INDIRECTREPLY_A_LOW_BITS] indirectreply_a_low_reg;
    reg      [`REG_INDIRECTREPLY_B_HI_BITS] indirectreply_b_hi_reg;
    reg      [`REG_INDIRECTREPLY_B_LOW_BITS] indirectreply_b_low_reg;
    reg      [`REG_INDIRECTCONFIG_BITS] indirectconfig_reg;
    reg      [`REG_INDIRECTCOMMAND_BITS] indirectcommand_reg;
    reg      [`REG_INDIRECTCOMMAND_BITS] indirectcommand_reg_internal;
    reg      indirectcommand_reg_update;

    // I/O Connections assignments
    assign S_AXI_AWREADY    = axi_awready;
    assign S_AXI_WREADY     = axi_wready;
    assign S_AXI_BRESP      = axi_bresp;
    assign S_AXI_BVALID     = axi_bvalid;
    assign S_AXI_ARREADY    = axi_arready;
    assign S_AXI_RDATA      = axi_rdata;
    assign S_AXI_RRESP      = axi_rresp;
    assign S_AXI_RVALID     = axi_rvalid;


    //Sample reset (not mandatory, but good practice)
    always @ (posedge clk) begin
        if (~resetn) begin
            resetn_sync_d  <=  1'b0;
            resetn_sync    <=  1'b0;
        end
        else begin
            resetn_sync_d  <=  resetn;
            resetn_sync    <=  resetn_sync_d;
        end
    end


    //global registers, sampling
    always @(posedge clk) resetn_soft <= #1 cpu_resetn_soft;

    // Implement axi_awready generation

    always @( posedge S_AXI_ACLK )
    begin
      if ( S_AXI_ARESETN == 1'b0 )
        begin
          axi_awready <= 1'b0;
        end
      else
        begin
          if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID)
            begin
              // slave is ready to accept write address when
              // there is a valid write address and write data
              // on the write address and data bus. This design
              // expects no outstanding transactions.
              axi_awready <= 1'b1;
            end
          else
            begin
              axi_awready <= 1'b0;
            end
        end
    end

    // Implement axi_awaddr latching

    always @( posedge S_AXI_ACLK )
    begin
      if ( S_AXI_ARESETN == 1'b0 )
        begin
          axi_awaddr <= 0;
        end
      else
        begin
          if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID)
            begin
              // Write Address latching
              axi_awaddr <= S_AXI_AWADDR ^ C_BASE_ADDRESS;
            end
        end
    end

    // Implement axi_wready generation

    always @( posedge S_AXI_ACLK )
    begin
      if ( S_AXI_ARESETN == 1'b0 )
        begin
          axi_wready <= 1'b0;
        end
      else
        begin
          if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID)
            begin
              // slave is ready to accept write data when
              // there is a valid write address and write data
              // on the write address and data bus. This design
              // expects no outstanding transactions.
              axi_wready <= 1'b1;
            end
          else
            begin
              axi_wready <= 1'b0;
            end
        end
    end

    // Implement write response logic generation

    always @( posedge S_AXI_ACLK )
    begin
      if ( S_AXI_ARESETN == 1'b0 )
        begin
          axi_bvalid  <= 0;
          axi_bresp   <= 2'b0;
        end
      else
        begin
          if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID)
            begin
              // indicates a valid write response is available
              axi_bvalid <= 1'b1;
              axi_bresp  <= 2'b0; // OKAY response
            end                   // work error responses in future
          else
            begin
              if (S_AXI_BREADY && axi_bvalid)
                //check if bready is asserted while bvalid is high)
                //(there is a possibility that bready is always asserted high)
                begin
                  axi_bvalid <= 1'b0;
                end
            end
        end
    end

    // Implement axi_arready generation

    always @( posedge S_AXI_ACLK )
    begin
      if ( S_AXI_ARESETN == 1'b0 )
        begin
          axi_arready <= 1'b0;
          axi_araddr  <= 32'b0;
        end
      else
        begin
          if (~axi_arready && S_AXI_ARVALID)
            begin
              // indicates that the slave has acceped the valid read address
              // Read address latching
              axi_arready <= 1'b1;
              axi_araddr  <= S_AXI_ARADDR ^ C_BASE_ADDRESS;
            end
          else
            begin
              axi_arready <= 1'b0;
            end
        end
    end


    // Implement axi_rvalid generation

    always @( posedge S_AXI_ACLK )
    begin
      if ( S_AXI_ARESETN == 1'b0 )
        begin
          axi_rvalid <= 0;
          axi_rresp  <= 0;
        end
      else
        begin
          if (axi_arready && S_AXI_ARVALID && ~axi_rvalid)
            begin
              // Valid read data is available at the read data bus
              axi_rvalid <= 1'b1;
              axi_rresp  <= 2'b0; // OKAY response
            end
          else if (axi_rvalid && S_AXI_RREADY)
            begin
              // Read data is accepted by the master
              axi_rvalid <= 1'b0;
            end
        end
    end


    // Implement memory mapped register select and write logic generation

    assign reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;

//////////////////////////////////////////////////////////////
// write registers
//////////////////////////////////////////////////////////////


//Write only register, clear on write (i.e. event)
    always @(posedge clk) begin
        if (!resetn_sync) begin
            reset_reg <= #1 `REG_RESET_DEFAULT;
        end
        else begin
            if (reg_wren) begin
                case (axi_awaddr)
                    //Reset Register
                        `REG_RESET_ADDR : begin
                                for ( byte_index = 0; byte_index <= (`REG_RESET_WIDTH/8-1); byte_index = byte_index +1)
                                    if (S_AXI_WSTRB[byte_index] == 1) begin
                                        reset_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8];
                                    end
                        end
                endcase
            end
            else begin
                reset_reg <= #1 `REG_RESET_DEFAULT;
            end
        end
    end

//R/W register, not cleared
    always @(posedge clk) begin
        if (!resetn_sync) begin

            cpu2ip_flip_reg <= #1 `REG_FLIP_DEFAULT;
            cpu2ip_debug_reg <= #1 `REG_DEBUG_DEFAULT;
            mac_0_hi_reg <= #1 `REG_MAC_0_HI_DEFAULT;
            mac_0_low_reg <= #1 `REG_MAC_0_LOW_DEFAULT;
            mac_1_hi_reg <= #1 `REG_MAC_1_HI_DEFAULT;
            mac_1_low_reg <= #1 `REG_MAC_1_LOW_DEFAULT;
            mac_2_hi_reg <= #1 `REG_MAC_2_HI_DEFAULT;
            mac_2_low_reg <= #1 `REG_MAC_2_LOW_DEFAULT;
            mac_3_hi_reg <= #1 `REG_MAC_3_HI_DEFAULT;
            mac_3_low_reg <= #1 `REG_MAC_3_LOW_DEFAULT;
            indirectaddress_reg <= #1 `REG_INDIRECTADDRESS_DEFAULT;
            indirectwrdata_a_hi_reg <= #1 `REG_INDIRECTREPLY_A_HI_DEFAULT;
            indirectwrdata_a_low_reg <= #1 `REG_INDIRECTREPLY_A_LOW_DEFAULT;
            indirectwrdata_b_hi_reg <= #1 `REG_INDIRECTREPLY_B_HI_DEFAULT;
            indirectwrdata_b_low_reg <= #1 `REG_INDIRECTREPLY_B_LOW_DEFAULT;
            indirectcommand_reg_internal <= #1 `REG_INDIRECTCOMMAND_DEFAULT;
            indirectconfig_reg <= #1 `REG_INDIRECTCONFIG_DEFAULT;
        end
        else begin
           if (reg_wren) //write event
            case (axi_awaddr)
            //Flip Register
                `REG_FLIP_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_FLIP_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            cpu2ip_flip_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //dynamic register;
                        end
                end
            //Debug Register
                `REG_DEBUG_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_DEBUG_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            cpu2ip_debug_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //dynamic register;
                        end
                end
            //Mac_0_hi Register
                `REG_MAC_0_HI_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_MAC_0_HI_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            mac_0_hi_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Mac_0_low Register
                `REG_MAC_0_LOW_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_MAC_0_LOW_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            mac_0_low_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Mac_1_hi Register
                `REG_MAC_1_HI_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_MAC_1_HI_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            mac_1_hi_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Mac_1_low Register
                `REG_MAC_1_LOW_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_MAC_1_LOW_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            mac_1_low_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Mac_2_hi Register
                `REG_MAC_2_HI_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_MAC_2_HI_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            mac_2_hi_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Mac_2_low Register
                `REG_MAC_2_LOW_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_MAC_2_LOW_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            mac_2_low_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Mac_3_hi Register
                `REG_MAC_3_HI_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_MAC_3_HI_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            mac_3_hi_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Mac_3_low Register
                `REG_MAC_3_LOW_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_MAC_3_LOW_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            mac_3_low_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Indirectaddress Register
                `REG_INDIRECTADDRESS_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_INDIRECTADDRESS_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            indirectaddress_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Indirectwrdata_a_hi Register
                `REG_INDIRECTWRDATA_A_HI_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_INDIRECTWRDATA_A_HI_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            indirectwrdata_a_hi_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Indirectwrdata_a_low Register
                `REG_INDIRECTWRDATA_A_LOW_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_INDIRECTWRDATA_A_LOW_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            indirectwrdata_a_low_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Indirectwrdata_b_hi Register
                `REG_INDIRECTWRDATA_B_HI_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_INDIRECTWRDATA_B_HI_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            indirectwrdata_b_hi_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Indirectwrdata_b_low Register
                `REG_INDIRECTWRDATA_B_LOW_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_INDIRECTWRDATA_B_LOW_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            indirectwrdata_b_low_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Indirectcommand Register
                `REG_INDIRECTCOMMAND_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_INDIRECTCOMMAND_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            indirectcommand_reg_internal[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
            //Indirectconfig Register         $finish;

                `REG_INDIRECTCONFIG_ADDR : begin
                    for ( byte_index = 0; byte_index <= (`REG_INDIRECTCONFIG_WIDTH/8-1); byte_index = byte_index +1)
                        if (S_AXI_WSTRB[byte_index] == 1) begin
                            indirectconfig_reg[byte_index*8 +: 8] <=  S_AXI_WDATA[byte_index*8 +: 8]; //static register;
                        end
                end
                default: begin
                end

            endcase
        end
   indirectcommand_reg_update <= reg_wren && (axi_awaddr == `REG_INDIRECTCOMMAND_ADDR);
  end



/////////////////////////
//// end of write
/////////////////////////

    // Implement memory mapped register select and read logic generation
    // Slave register read enable is asserted when valid address is available
    // and the slave is ready to accept the read address.

    // reg_rden control logic
    // temperary no extra logic here
    assign reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;

    always @(*)
    begin

        case ( axi_araddr /*S_AXI_ARADDR ^ C_BASE_ADDRESS*/)
            //Id Register
            `REG_ID_ADDR : begin
                reg_data_out [`REG_ID_BITS] =  id_reg;
            end
            //Version Register
            `REG_VERSION_ADDR : begin
                reg_data_out [`REG_VERSION_BITS] =  version_reg;
            end
            //Flip Register
            `REG_FLIP_ADDR : begin
                reg_data_out [`REG_FLIP_BITS] =  ip2cpu_flip_reg;
            end
            //Debug Register
            `REG_DEBUG_ADDR : begin
                reg_data_out [`REG_DEBUG_BITS] =  ip2cpu_debug_reg;
            end
            //Pkt_sent_from_cpu_cntr Register
            `REG_PKT_SENT_FROM_CPU_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_SENT_FROM_CPU_CNTR_BITS] =  pkt_sent_from_cpu_cntr_reg;
            end
            //Pkt_sent_to_cpu_options_ver_cntr Register
            `REG_PKT_SENT_TO_CPU_OPTIONS_VER_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_SENT_TO_CPU_OPTIONS_VER_CNTR_BITS] =  pkt_sent_to_cpu_options_ver_cntr_reg;
            end
            //Pkt_sent_to_cpu_bad_ttl_cntr Register
            `REG_PKT_SENT_TO_CPU_BAD_TTL_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_SENT_TO_CPU_BAD_TTL_CNTR_BITS] =  pkt_sent_to_cpu_bad_ttl_cntr_reg;
            end
            //Pkt_sent_to_cpu_dest_ip_hit_cntr Register
            `REG_PKT_SENT_TO_CPU_DEST_IP_HIT_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_SENT_TO_CPU_DEST_IP_HIT_CNTR_BITS] =  pkt_sent_to_cpu_dest_ip_hit_cntr_reg;
            end
            //Pkt_forwarded_cntr Register
            `REG_PKT_FORWARDED_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_FORWARDED_CNTR_BITS] =  pkt_forwarded_cntr_reg;
            end
            //Pkt_dropped_checksum_cntr Register
            `REG_PKT_DROPPED_CHECKSUM_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_DROPPED_CHECKSUM_CNTR_BITS] =  pkt_dropped_checksum_cntr_reg;
            end
            //Pkt_sent_to_cpu_non_ip_cntr Register
            `REG_PKT_SENT_TO_CPU_NON_IP_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_SENT_TO_CPU_NON_IP_CNTR_BITS] =  pkt_sent_to_cpu_non_ip_cntr_reg;
            end
            //Pkt_sent_to_cpu_arp_miss_cntr Register
            `REG_PKT_SENT_TO_CPU_ARP_MISS_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_SENT_TO_CPU_ARP_MISS_CNTR_BITS] =  pkt_sent_to_cpu_arp_miss_cntr_reg;
            end
            //Pkt_sent_to_cpu_lpm_miss_cntr Register
            `REG_PKT_SENT_TO_CPU_LPM_MISS_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_SENT_TO_CPU_LPM_MISS_CNTR_BITS] =  pkt_sent_to_cpu_lpm_miss_cntr_reg;
            end
            //Pkt_dropped_wrong_dst_mac_cntr Register
            `REG_PKT_DROPPED_WRONG_DST_MAC_CNTR_ADDR : begin
                reg_data_out [`REG_PKT_DROPPED_WRONG_DST_MAC_CNTR_BITS] =  pkt_dropped_wrong_dst_mac_cntr_reg;
            end
            //Mac_0_hi Register
            `REG_MAC_0_HI_ADDR : begin
                reg_data_out [`REG_MAC_0_HI_BITS] =  mac_0_hi_reg;
            end
            //Mac_0_low Register
            `REG_MAC_0_LOW_ADDR : begin
                reg_data_out [`REG_MAC_0_LOW_BITS] =  mac_0_low_reg;
            end
            //Mac_1_hi Register
            `REG_MAC_1_HI_ADDR : begin
                reg_data_out [`REG_MAC_1_HI_BITS] =  mac_1_hi_reg;
            end
            //Mac_1_low Register
            `REG_MAC_1_LOW_ADDR : begin
                reg_data_out [`REG_MAC_1_LOW_BITS] =  mac_1_low_reg;
            end
            //Mac_2_hi Register
            `REG_MAC_2_HI_ADDR : begin
                reg_data_out [`REG_MAC_2_HI_BITS] =  mac_2_hi_reg;
            end
            //Mac_2_low Register
            `REG_MAC_2_LOW_ADDR : begin
                reg_data_out [`REG_MAC_2_LOW_BITS] =  mac_2_low_reg;
            end
            //Mac_3_hi Register
            `REG_MAC_3_HI_ADDR : begin
                reg_data_out [`REG_MAC_3_HI_BITS] =  mac_3_hi_reg;
            end
            //Mac_3_low Register
            `REG_MAC_3_LOW_ADDR : begin
                reg_data_out [`REG_MAC_3_LOW_BITS] =  mac_3_low_reg;
	    end
            //Indirectaddress Register
            `REG_INDIRECTADDRESS_ADDR : begin
                reg_data_out [`REG_INDIRECTADDRESS_BITS] =  indirectaddress_reg;
            end
            //Indirectwrdata_a_hi Register
            `REG_INDIRECTWRDATA_A_HI_ADDR : begin
                reg_data_out [`REG_INDIRECTWRDATA_A_HI_BITS] =  indirectwrdata_a_hi_reg;
            end
            //Indirectwrdata_a_low Register
            `REG_INDIRECTWRDATA_A_LOW_ADDR : begin
                reg_data_out [`REG_INDIRECTWRDATA_A_LOW_BITS] =  indirectwrdata_a_low_reg;
            end
            //Indirectwrdata_b_hi Register
            `REG_INDIRECTWRDATA_B_HI_ADDR : begin
                reg_data_out [`REG_INDIRECTWRDATA_B_HI_BITS] =  indirectwrdata_b_hi_reg;
            end
            //Indirectwrdata_b_low Register
            `REG_INDIRECTWRDATA_B_LOW_ADDR : begin
                reg_data_out [`REG_INDIRECTWRDATA_B_LOW_BITS] =  indirectwrdata_b_low_reg;
            end
            //Indirectreply_a_hi Register
            `REG_INDIRECTREPLY_A_HI_ADDR : begin
                reg_data_out [`REG_INDIRECTREPLY_A_HI_BITS] =  indirectreply_a_hi_reg;
            end
            //Indirectreply_a_low Register
            `REG_INDIRECTREPLY_A_LOW_ADDR : begin
                reg_data_out [`REG_INDIRECTREPLY_A_LOW_BITS] =  indirectreply_a_low_reg;
            end
            //Indirectreply_b_hi Register
            `REG_INDIRECTREPLY_B_HI_ADDR : begin
                reg_data_out [`REG_INDIRECTREPLY_B_HI_BITS] =  indirectreply_b_hi_reg;
            end
            //Indirectreply_b_low Register
            `REG_INDIRECTREPLY_B_LOW_ADDR : begin
                reg_data_out [`REG_INDIRECTREPLY_B_LOW_BITS] =  indirectreply_b_low_reg;
            end
            //Indirectcommand Register
            `REG_INDIRECTCOMMAND_ADDR : begin
                reg_data_out [`REG_INDIRECTCOMMAND_BITS] =  indirectcommand_reg;
            end
            //Indirectconfig Register
            `REG_INDIRECTCONFIG_ADDR : begin
                reg_data_out [`REG_INDIRECTCONFIG_BITS] =  indirectconfig_reg;
            end
            //Default return value
            default: begin
                reg_data_out [31:0] =  32'hDEADBEEF;
            end

        endcase

    end//end of assigning data to IP2Bus_Data bus

    //Read only registers, not cleared
    //Nothing to do here....

//Read only registers, cleared on read (e.g. counters)
    always @(posedge clk)
    if (!resetn_sync) begin
        pkt_sent_from_cpu_cntr_reg_clear <= #1 1'b0;
        pkt_sent_from_cpu_cntr_reg_clear_d <= #1 1'b0;
        pkt_sent_to_cpu_options_ver_cntr_reg_clear <= #1 1'b0;
        pkt_sent_to_cpu_options_ver_cntr_reg_clear_d <= #1 1'b0;
        pkt_sent_to_cpu_bad_ttl_cntr_reg_clear <= #1 1'b0;
        pkt_sent_to_cpu_bad_ttl_cntr_reg_clear_d <= #1 1'b0;
        pkt_sent_to_cpu_dest_ip_hit_cntr_reg_clear <= #1 1'b0;
        pkt_sent_to_cpu_dest_ip_hit_cntr_reg_clear_d <= #1 1'b0;
        pkt_forwarded_cntr_reg_clear <= #1 1'b0;
        pkt_forwarded_cntr_reg_clear_d <= #1 1'b0;
        pkt_dropped_checksum_cntr_reg_clear <= #1 1'b0;
        pkt_dropped_checksum_cntr_reg_clear_d <= #1 1'b0;
        pkt_sent_to_cpu_non_ip_cntr_reg_clear <= #1 1'b0;
        pkt_sent_to_cpu_non_ip_cntr_reg_clear_d <= #1 1'b0;
        pkt_sent_to_cpu_arp_miss_cntr_reg_clear <= #1 1'b0;
        pkt_sent_to_cpu_arp_miss_cntr_reg_clear_d <= #1 1'b0;
        pkt_sent_to_cpu_lpm_miss_cntr_reg_clear <= #1 1'b0;
        pkt_sent_to_cpu_lpm_miss_cntr_reg_clear_d <= #1 1'b0;
        pkt_dropped_wrong_dst_mac_cntr_reg_clear <= #1 1'b0;
        pkt_dropped_wrong_dst_mac_cntr_reg_clear_d <= #1 1'b0;
    end
    else begin
        pkt_sent_from_cpu_cntr_reg_clear <= #1 pkt_sent_from_cpu_cntr_reg_clear_d;
        pkt_sent_from_cpu_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_SENT_FROM_CPU_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_sent_to_cpu_options_ver_cntr_reg_clear <= #1 pkt_sent_to_cpu_options_ver_cntr_reg_clear_d;
        pkt_sent_to_cpu_options_ver_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_SENT_TO_CPU_OPTIONS_VER_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_sent_to_cpu_bad_ttl_cntr_reg_clear <= #1 pkt_sent_to_cpu_bad_ttl_cntr_reg_clear_d;
        pkt_sent_to_cpu_bad_ttl_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_SENT_TO_CPU_BAD_TTL_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_sent_to_cpu_dest_ip_hit_cntr_reg_clear <= #1 pkt_sent_to_cpu_dest_ip_hit_cntr_reg_clear_d;
        pkt_sent_to_cpu_dest_ip_hit_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_SENT_TO_CPU_DEST_IP_HIT_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_forwarded_cntr_reg_clear <= #1 pkt_forwarded_cntr_reg_clear_d;
        pkt_forwarded_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_FORWARDED_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_dropped_checksum_cntr_reg_clear <= #1 pkt_dropped_checksum_cntr_reg_clear_d;
        pkt_dropped_checksum_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_DROPPED_CHECKSUM_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_sent_to_cpu_non_ip_cntr_reg_clear <= #1 pkt_sent_to_cpu_non_ip_cntr_reg_clear_d;
        pkt_sent_to_cpu_non_ip_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_SENT_TO_CPU_NON_IP_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_sent_to_cpu_arp_miss_cntr_reg_clear <= #1 pkt_sent_to_cpu_arp_miss_cntr_reg_clear_d;
        pkt_sent_to_cpu_arp_miss_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_SENT_TO_CPU_ARP_MISS_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_sent_to_cpu_lpm_miss_cntr_reg_clear <= #1 pkt_sent_to_cpu_lpm_miss_cntr_reg_clear_d;
        pkt_sent_to_cpu_lpm_miss_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_SENT_TO_CPU_LPM_MISS_CNTR_ADDR)) ? 1'b1 : 1'b0;
        pkt_dropped_wrong_dst_mac_cntr_reg_clear <= #1 pkt_dropped_wrong_dst_mac_cntr_reg_clear_d;
        pkt_dropped_wrong_dst_mac_cntr_reg_clear_d <= #1(reg_rden && (axi_araddr==`REG_PKT_DROPPED_WRONG_DST_MAC_CNTR_ADDR)) ? 1'b1 : 1'b0;
    end


// Output register or memory read data
    always @( posedge S_AXI_ACLK )
    begin
      if ( S_AXI_ARESETN == 1'b0 )
        begin
          axi_rdata  <= 0;
        end
      else
        begin
          // When there is a valid read address (S_AXI_ARVALID) with
          // acceptance of read address by the slave (axi_arready),
          // output the read dada
          if (reg_rden)
            begin
              axi_rdata <= reg_data_out/*ip2bus_data*/;     // register read data /* some new changes here */
            end
        end
    end

    //////////////////////////////////
    // Implement Indirect Access
	//////////////////////////////////
	

  //--------------------- Internal Parameters-------------------------
   localparam NUM_INDIRECT_STATES                = 6;
   localparam IDLE_INDIRECT_STATE                = 1;
   localparam WRITE_INDIRECT_STATE               = 2;
   localparam WRITE_WAIT_INDIRECT_STATE          = 4;
   localparam READ_INDIRECT_STATE                = 8;
   localparam READ_WAIT_INDIRECT_STATE           = 16;
   localparam INDIRECT_DONE_STATE                = 32;
   localparam INDIRECT_WRITE                     = 0;
   localparam INDIRECT_READ                      = 1;
   localparam INDIRECT_WRITE_TA                  = 1;
   localparam INDIRECT_WRITE_WS                  = 0;
  //------------------------------------------------------------------
   
   reg  [NUM_INDIRECT_STATES-1:0]           indirect_state, indirect_state_next, indirect_state_last;
   wire                            indirect_trigger;
   wire                            indirect_type;
   reg                             indirect_status, indirect_status_next;
   wire [3:0]                      indirect_address_increment;
   wire                            indirect_write_type;
   wire [10:0]                     indirect_timeout;
   wire [15:0]                     indirect_repeat_count;
   reg  [15:0]                     indirect_remaining,indirect_remaining_next;
   reg  [10:0]                     indirect_timeout_count, indirect_timeout_count_next;
   reg                             indirect_reply_valid;
   reg  [31:0]                     indirect_address,indirect_address_next;
   reg  [3:0]                      indirect_memory_select,indirect_memory_select_next;
   wire                             indirect_command_done;
   
   assign   indirect_trigger = indirectcommand_reg[0];
   assign   indirect_type    = indirectcommand_reg[4];
   assign   indirect_address_increment = indirectconfig_reg[3:0];
   assign   indirect_write_type = indirectconfig_reg[4];
   assign   indirect_timeout    = indirectconfig_reg[15:5];
   assign   indirect_repeat_count = indirectconfig_reg[31:16];
   
 always @(*) begin
      indirect_state_next   = indirect_state;
      indirect_status_next  = indirect_status;
      indirect_remaining_next = indirect_remaining;
      indirect_timeout_count_next = indirect_timeout_count;
      indirect_address_next      = indirect_address;
      indirect_memory_select_next = indirect_memory_select;
      case(indirect_state)
        IDLE_INDIRECT_STATE: begin
     	   if(indirect_trigger) begin
     	      indirect_state_next= (indirect_type == INDIRECT_WRITE) ? WRITE_INDIRECT_STATE : READ_INDIRECT_STATE;
     	      indirect_remaining_next = (indirect_repeat_count == 0) ? 16'h1 : indirect_repeat_count;
     	      indirect_timeout_count_next   = indirect_timeout;
     	      indirect_address_next   =  indirectaddress_reg; //This is the address in the user register
     	      indirect_memory_select_next = indirectaddress_reg[31:28];
     	   end
	    end
	    
	    READ_INDIRECT_STATE: begin
		     indirect_state_next = READ_WAIT_INDIRECT_STATE;
	    end
	    READ_WAIT_INDIRECT_STATE: begin
	         if (indirect_reply_valid) begin
	            indirect_state_next = INDIRECT_DONE_STATE;
	            indirect_status_next =0;
	         end
	         if (indirect_timeout_count==0) begin
	            indirect_state_next = INDIRECT_DONE_STATE;
	            indirect_status_next = 1; 
	         end
	         indirect_timeout_count_next = indirect_timeout_count-1;
	     end
	     WRITE_INDIRECT_STATE: begin
	         indirect_state_next = WRITE_WAIT_INDIRECT_STATE;
	     end
	     WRITE_WAIT_INDIRECT_STATE:  begin
	         if (((indirect_write_type == INDIRECT_WRITE_TA) && (indirect_reply_valid)) || ((indirect_write_type == INDIRECT_WRITE_WS) && (indirect_timeout_count==0))) begin
	           indirect_remaining_next = indirect_remaining - 1;
	           indirect_address_next = indirect_address+indirect_address_increment;
	           if (indirect_remaining==1) begin
	              indirect_state_next = INDIRECT_DONE_STATE;
	           end
	         end
	         else 
	           if (indirect_timeout_count==0) begin
	         	indirect_state_next = INDIRECT_DONE_STATE;
	         	indirect_status_next = 1; 
	         end
             indirect_timeout_count_next = indirect_timeout_count==0 ? 0 : indirect_timeout_count-1;
	     end
	     INDIRECT_DONE_STATE: begin
	        indirect_state_next= IDLE_INDIRECT_STATE;
	     end
	     default: begin
	         indirect_state_next= IDLE_INDIRECT_STATE;
	     end
      endcase // case(state)
   end // always @ (*)
   
    assign indirect_command_done = (indirect_state==INDIRECT_DONE_STATE);
   
   always @(posedge clk) begin
      if(~resetn_sync) begin
         indirect_state <= #1 IDLE_INDIRECT_STATE;
         indirect_state_last <= #1 IDLE_INDIRECT_STATE;
         indirect_status <= #1 1'b0;
         indirect_remaining <= #1 0;
         indirect_timeout_count <= #1 0;
         indirect_address   <= #1 0;
         indirect_memory_select <= #1 0;
         indirectcommand_reg <= #1 `REG_INDIRECTCOMMAND_DEFAULT;
      end
      else begin
         indirect_state <= #1 indirect_state_next;
         indirect_state_last <= #1 indirect_state;
         indirect_status <= #1 indirect_status_next;
         indirect_remaining <= #1 indirect_remaining_next;
         indirect_timeout_count <= #1 indirect_timeout_count_next;
         indirect_address   <= #1  indirect_address_next;
         indirect_memory_select <= #1 indirect_memory_select_next;
         indirectcommand_reg <= #1  indirect_command_done ? {indirect_status,indirectcommand_reg[7:4],4'h0} : 
                                    indirectcommand_reg_update ? indirectcommand_reg_internal: 
                                    indirectcommand_reg;
      end
   end   
   

       
       always @(posedge clk) begin
         if  (~resetn_sync) begin
           ip_lpm_tcam_addr <= #1 0;
           ip_lpm_tcam_data <= #1 0;
           ip_lpm_tcam_rd_wrn<= #1 0;
           ip_lpm_tcam_cmd_valid <= #1 0;
         end 
         else begin
           ip_lpm_tcam_addr <= #1 indirect_address;
           ip_lpm_tcam_data <= #1 {indirectwrdata_a_hi_reg,indirectwrdata_a_low_reg,indirectwrdata_b_hi_reg,indirectwrdata_b_low_reg};
           ip_lpm_tcam_rd_wrn<= #1 indirect_type;
           ip_lpm_tcam_cmd_valid <= #1 (32'h00000000==(indirect_memory_select<<28)) && ((indirect_state == WRITE_INDIRECT_STATE) || (indirect_state == READ_INDIRECT_STATE));
         end 
       end

       
       always @(posedge clk) begin
         if  (~resetn_sync) begin
           ip_arp_cam_addr <= #1 0;
           ip_arp_cam_data <= #1 0;
           ip_arp_cam_rd_wrn<= #1 0;
           ip_arp_cam_cmd_valid <= #1 0;
         end 
         else begin
           ip_arp_cam_addr <= #1 indirect_address;
           ip_arp_cam_data <= #1 {indirectwrdata_a_hi_reg,indirectwrdata_a_low_reg,indirectwrdata_b_hi_reg,indirectwrdata_b_low_reg};
           ip_arp_cam_rd_wrn<= #1 indirect_type;
           ip_arp_cam_cmd_valid <= #1 (32'h10000000==(indirect_memory_select<<28)) && ((indirect_state == WRITE_INDIRECT_STATE) || (indirect_state == READ_INDIRECT_STATE));
         end 
       end

       
       always @(posedge clk) begin
         if  (~resetn_sync) begin
           dest_ip_cam_addr <= #1 0;
           dest_ip_cam_data <= #1 0;
           dest_ip_cam_rd_wrn<= #1 0;
           dest_ip_cam_cmd_valid <= #1 0;
         end 
         else begin
           dest_ip_cam_addr <= #1 indirect_address;
           dest_ip_cam_data <= #1 {indirectwrdata_a_hi_reg,indirectwrdata_a_low_reg,indirectwrdata_b_hi_reg,indirectwrdata_b_low_reg};
           dest_ip_cam_rd_wrn<= #1 indirect_type;
           dest_ip_cam_cmd_valid <= #1 (32'h20000000==(indirect_memory_select<<28)) && ((indirect_state == WRITE_INDIRECT_STATE) || (indirect_state == READ_INDIRECT_STATE));
         end 
       end

       always @(posedge clk) begin
          if  (~resetn_sync) begin
             indirectreply_a_hi_reg <= #1 0;
             indirectreply_a_low_reg <= #1 0;
             indirectreply_b_hi_reg <= #1 0;
             indirectreply_b_low_reg <= #1 0;
             indirect_reply_valid <= #1 0; 
          end 
          else begin 
             indirectreply_a_hi_reg <= #1 32'h00000000==(indirect_memory_select<<28) ? ip_lpm_tcam_reply[127:96] :32'h10000000==(indirect_memory_select<<28) ? ip_arp_cam_reply[127:96] :32'h20000000==(indirect_memory_select<<28) ? dest_ip_cam_reply[127:96] : 0;
            indirectreply_a_low_reg <= #1 32'h00000000==(indirect_memory_select<<28) ? ip_lpm_tcam_reply[95:64] :32'h10000000==(indirect_memory_select<<28) ? ip_arp_cam_reply[95:64] :32'h20000000==(indirect_memory_select<<28) ? dest_ip_cam_reply[95:64] : 0;
             indirectreply_b_hi_reg <= #1 32'h00000000==(indirect_memory_select<<28) ? ip_lpm_tcam_reply[63:32] :32'h10000000==(indirect_memory_select<<28) ? ip_arp_cam_reply[63:32] :32'h20000000==(indirect_memory_select<<28) ? dest_ip_cam_reply[63:32] : 0;
             indirectreply_b_low_reg <= #1 32'h00000000==(indirect_memory_select<<28) ? ip_lpm_tcam_reply[31:0] :32'h10000000==(indirect_memory_select<<28) ? ip_arp_cam_reply[31:0] :32'h20000000==(indirect_memory_select<<28) ? dest_ip_cam_reply[31:0] : 0;
             indirect_reply_valid <= #1 32'h00000000==(indirect_memory_select<<28) ? ip_lpm_tcam_reply_valid :32'h10000000==(indirect_memory_select<<28) ? ip_arp_cam_reply_valid :32'h20000000==(indirect_memory_select<<28) ? dest_ip_cam_reply_valid : 0;
          end 
        end
  
endmodule
